`ifndef _PARAMETER_VH_
`define _PARAMETER_VH_

`define DECLARE_MODE_PARAMETERS \
    localparam TRAIN = 1'b1, \
               TEST  = 1'b0;

`endif
