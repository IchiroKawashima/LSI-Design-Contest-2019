`ifndef _PARAMETER_VH_
`define _PARAMETER_VH_

// Number of Neurons
`define PARAM_NB_INPUT_NEURON 100
`define PARAM_NB_HIDDEN0_NEURON 100
`define PARAM_NB_HIDDEN1_NEURON 100
`define PARAM_NB_OUTPUT_NEURON 100

// Bit Width
`define PARAM_SYNAPSE_BITWIDTH 8
`define PARAM_NEURON_BITWIDTH 8

`define DECLARE_PARAMETERS \
    localparam NB_INPUT_NEURON   = `PARAM_NB_INPUT_NEURON; \
    localparam NB_HIDDEN0_NEURON = `PARAM_NB_HIDDEN0_NEURON; \
    localparam NB_HIDDEN1_NEURON = `PARAM_NB_HIDDEN1_NEURON; \
    localparam NB_OUTPUT_NEURON  = `PARAM_NB_OUTPUT_NEURON; \
    localparam SYNAPSE_BITWIDTH  = `PARAM_SYNAPSE_BITWIDTH; \
    localparam NEURON_BITWIDTH   = `PARAM_NEURON_BITWIDTH;

`endif
